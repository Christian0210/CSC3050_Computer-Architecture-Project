`timescale 1ns/1ps

module alu_test;

reg[31:0] i_datain,gr1,gr2;
reg[31:0] imm;

wire[31:0] c;
wire zero;
wire overflow;
wire neg;

alu testalu(i_datain,gr1,gr2,c,imm,zero,neg,overflow);

initial
begin
    // add func:00 op:00
    $display("\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SLL TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    $monitor("   %h : %h :  %h  |%h:%h:%h:%h|%h:%h:%h:%h|  %h   :  %h  :   %h",
    i_datain, testalu.opcode, testalu.func, gr1, gr2, c, imm, testalu.reg_A, testalu.reg_B, testalu.reg_C, testalu.Imm, zero, neg, overflow);
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0000;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_1000_0000;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0000;
    gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0001_0000_0000;
    gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    #10

    // sllv func: 02 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SRL TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0010;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_1000_0010;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0010;
    gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0001_0000_0010;
    gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    #10

    // sllv func: 03 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SRA TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0011;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_1000_0011;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0100_0011;
    gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0001_0000_0011;
    gr2<=32'b0100_0000_0100_0000_0100_0000_0100_0000;
    #10

    // sllv func: 04 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SLLV TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0100;
    gr1<=32'b1;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0100;
    gr1<=32'b10;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10

    // srlv func: 06 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SRLV TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0110;
    gr1<=32'b1;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0110;
    gr1<=32'b10;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10
    
    // srav func: 07 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SRAV TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0111;
    gr1<=32'b1;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0000_0111;
    gr1<=32'b10;
    gr2<=32'b1101_1101_1101_1101_1101_1101_1101_1101;
    #10

     // add func: 18 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_MULT TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1000;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1000;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10


    // add func: 19 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_MULTU TEST                                                  ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1001;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1001;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10


    // add func: 1a op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_DIV TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1010;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1010;
    //gr1     <=32'b1000_0000_0000_0000_0000_0000_0001_0001;
    gr1     <=32'b1111_1111_1111_1111_1111_1111_1110_1111;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10


    // add func: 1b op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_DIVU TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1011;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0001_1011;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10

    // add func: 20 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_ADD TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
    gr1     <=32'b1010_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b1011_1111_1111_1111_1111_1111_1111_1111;//negative overflow
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
    gr1     <=32'b0111_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b0111_1111_1001_1111_0001_1111_1111_1111;//positive overflow
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000;
    gr1     <=32'b1111_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b10;//negative flag
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0000; 
    gr1     <=32'b0;
    gr2     <=32'b0;//zero
    #10

    // add func: 21 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_ADDU TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
    gr1     <=32'b1010_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b1011_1111_1111_1111_1111_1111_1111_1111;//no negative overflow
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
    gr1     <=32'b0111_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b0111_1111_1001_1111_0001_1111_1111_1111;//no positive overflow
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001;
    gr1     <=32'b1111_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b10;//negative flag
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0001; 
    gr1     <=32'b0;
    gr2     <=32'b0;//zero
    #10

    // add func: 22 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SUB TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
    gr1     <=32'b10;
    gr2     <=32'b1100;//negative flag
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
    gr1     <=32'b0111_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b1011_1111_1111_1111_1111_1111_1111_1111;//negative overflow
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010; 
    gr1     <=32'b1011_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b0111_1111_1111_1111_1101_1111_1111_1111;//positive overflow
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0010;
    gr1     <=32'b0;
    gr2     <=32'b0;//zero
    #10

    // add func: 23 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SUBU TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
    gr1     <=32'b10;
    gr2     <=32'b1100;//negative flag
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
    gr1     <=32'b0111_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b1011_1111_1111_1111_1111_1111_1111_1111;//no negative overflow
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011; 
    gr1     <=32'b1011_1111_1111_1111_1111_1111_1111_1011;
    gr2     <=32'b0111_1111_1111_1111_1101_1111_1111_1111;//no positive overflow
    #10 
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0011;
    gr1     <=32'b0;
    gr2     <=32'b0;//zero
    #10

    // add func: 24 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_AND TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0100;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0001_0000_0001_0000;
    #10

    // xor func: 25 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_OR TEST                                                     ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0101;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0001_0000_0001_0000;
    #10

    // xor func: 26 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_XOR TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0110;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0001_0000_0001_0000;
    #10

    // add func: 27 op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_NOR TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_0111;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0001_0000_0001_0000;
    #10
  
    // slt func: 2a op: 00
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SLT TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b1000_0000_0000_0000_0000_0000_0000_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1010;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0000_0001;
    gr2     <=32'b1000_0000_0000_0000_0000_0000_0001_0001;
    #10

    // sltu func: 2b op: 00  
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SLTU TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b1000_0000_0000_0000_0000_0000_0000_0001;
    #10
    i_datain<=32'b0000_0000_0000_0001_0001_0000_0010_1011;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0000_0001;
    gr2     <=32'b1000_0000_0000_0000_0000_0000_0001_0001;
    #10

    // add op: 04
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_BEQ TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0001_0000_0000_0000_0000_0000_1111_1111;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0001_0000_0000_0000_0000_0000_1111_1111;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    #10

    // add op: 05
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_BNE TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0001_0100_0000_0000_0000_0000_1111_1111;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    #10
    i_datain<=32'b0001_0100_0000_0000_0000_0000_1111_1111;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0000_0000_0000_0001;
    #10

    // add op: 08
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_ADDI TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0010_0000_0000_0000_0000_0000_0001_0001;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0;
    #10
    i_datain<=32'b0010_0000_0000_0000_1000_0000_0001_0001;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0000_0001;//negative overflow
    gr2     <=32'b0;
    #10 
    i_datain<=32'b0010_0000_0000_0000_0000_0000_0001_0001;
    gr1     <=32'b0111_1111_1111_1111_1111_1111_1111_1111;//positive overflow
    gr2     <=32'b0;
    #10 
    i_datain<=32'b0010_0000_0000_0000_0000_0000_0001_0001;
    gr1     <=32'b1111_0000_0000_0000_0000_0000_0000_0001;//negative flag
    gr2     <=32'b0;
    #10
    i_datain<=32'b0010_0000_0000_0000_0000_0000_0000_0000;
    gr1     <=32'b0;//zero
    gr2     <=32'b0;
    #10

    // add op: 09
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_ADDIU TEST                                                  ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0010_0100_0000_0000_0000_0000_0001_0001;
    gr1     <=32'b0000_0000_0000_0000_0000_0000_0001_0001;
    gr2     <=32'b0;
    #10
    i_datain<=32'b0010_0100_0000_0000_1000_0000_0001_0001;
    gr1     <=32'b1000_0000_0000_0000_0000_0000_0000_0001;//no negative overflow
    gr2     <=32'b0;
    #10 
    i_datain<=32'b0010_0100_0000_0000_0000_0000_0001_0001;
    gr1     <=32'b0111_1111_1111_1111_1111_1111_1111_1111;//no positive overflow
    gr2     <=32'b0;
    #10 
    i_datain<=32'b0010_0100_0000_0000_0000_0000_0001_0001;
    gr1     <=32'b1111_0000_0000_0000_0000_0000_0000_0001;//negative flag
    gr2     <=32'b0;
    #10
    i_datain<=32'b0010_0100_0000_0000_0000_0000_0000_0000;
    gr1     <=32'b0;//zero
    gr2     <=32'b0;
    #10

    // add op: 0a
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SLTI TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0010_1000_0000_0000_0000_0001_0000_0001;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0;
    #10
    i_datain<=32'b0010_1000_0000_0000_0001_0001_0001_0001;
    gr1     <=32'b0000_0000_0000_0000_0000_0001_0000_0001;
    gr2     <=32'b0;
    #10

    // xor op: 0b
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SLTIU TEST                                                  ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0010_1100_0000_0000_0000_0001_0000_0001;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0;
    #10
    i_datain<=32'b0010_1100_0000_0000_0001_0001_0001_0001;
    gr1     <=32'b0000_0000_0000_0000_0000_0001_0000_0001;
    gr2     <=32'b0;
    #10


    // add op: 0c
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_ANDI TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0011_0000_0000_0000_0000_0001_0000_0001;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0000_0000_0000_0000_0001_0000_0001_0000;
    #10

    // xor op: 0d
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_ORI TEST                                                    ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0011_0100_0000_0000_0000_0001_0000_0001;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0;
    #10

    // xor op: 0e
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_XORI TEST                                                   ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b0011_1000_0000_0000_0000_0001_0000_0001;
    gr1     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    gr2     <=32'b0;
    #10

    // lw op: 23
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_LW TEST                                                     ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b1000_1100_0000_0000_0000_0000_1111_1111;
    gr1     <=32'b0;
    gr2     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;
    #10

    // sw op: 2b
    $display("\n\n");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("                                                     MIPS_SW TEST                                                     ");
    $display("----------------------------------------------------------------------------------------------------------------------");
    $display("      instruction       |                              parameter                                |         flag        ");
    $display("instruction : op : func |  gr1   :  gr2   :   c    :  imm   | reg_A  : reg_B  : reg_C  :  Imm   | zero : neg :overflow");
    i_datain<=32'b1010_1100_0000_0000_0000_0000_1111_1111;
    gr1     <=32'b0;
    gr2     <=32'b0000_0000_0000_0000_0001_0001_0001_0001;

    $finish;
end
endmodule